module core (
    
);
    
endmodule
    
endmodule